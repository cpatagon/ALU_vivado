lgomez@meteo.9542:1723388680
lgomez@meteo.77839:1723295069